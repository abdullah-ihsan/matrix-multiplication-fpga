module top (
    input wire clk,  // System clock
    input wire rst,  // Reset
    input wire rx,   // UART RX
    output wire tx   // UART TX
);
    // Instantiate UART RX/TX modules
    // Instantiate memory modules for matrices A, B, and C
    // Instantiate matrix multiplication module
    // Instantiate FSM for control
endmodule
